///// verilog code for xnor gate design

module xnor_gate( input a, b, output y);

xnor(y, a, b);

endmodule







