/// Verilog code for OR gate
module or_gate(input a, b, output y);

assign y = a | b;

endmodule
